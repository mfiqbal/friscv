module tester;
endmodule
