`ifndef FARM_PKG
`define FARM_PKG

package farm_pkg;
	`define cq 3  // clock to q delay
	`define cd 3  // combinational delay 
endpackage


`endif
